//============================================================================
//
//  Memory tester for MiSTer.              https://github.com/MiSTer-devel/MemTest_MiSTer
//  Copyright (C) 2017-2019 Sorgelig
//
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//
//  You should have received a copy of the GNU General Public License along
//  with this program; if not, write to the Free Software Foundation, Inc.,
//  51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.
//============================================================================
//============================================================================
//
//  Multicore 2 Top by Victor Trucco
//
//============================================================================
//============================================================================
//
//  neptUNO Top adapted by delgrom         https://github.com/neptuno-fpga/MemTest_Mister
//
//============================================================================
//============================================================================
//
//  DECA Top adapted by somhic
//
//============================================================================


`default_nettype none

module memtest_deca
( 
	// Clocks
	input wire	clock_50_i,

	// KEY / SW
	input 		     [1:0]		KEY,
	input 		     [1:0]		SW,
	
	// SDRAM	
	output [12:0] SDRAM_A,
	output  [1:0] SDRAM_BA,
	inout  [15:0] SDRAM_DQ,
	output        SDRAM_DQMH,
	output        SDRAM_DQML,
	output        SDRAM_CKE,
	output        SDRAM_nCS,
	output        SDRAM_nWE,
	output        SDRAM_nRAS,
	output        SDRAM_nCAS,
	output        SDRAM_CLK,

	// PS2
	input wire	ps2_clk_io,
	input wire	ps2_data_io,

        // Joysticks    
	/* output wire joy_clock_o       = 1'b1,
	   output wire joy_load_o        = 1'b1,
	   input  wire joy_data_i,
	   output wire joy_p7_o          = 1'b1,
        */

	// HDMI-TX 
	inout 		          		HDMI_I2C_SCL,
	inout 		          		HDMI_I2C_SDA,
	inout 		     [3:0]		HDMI_I2S,
	inout 		          		HDMI_LRCLK,
	inout 		          		HDMI_MCLK,
	inout 		          		HDMI_SCLK,
	output		          		HDMI_TX_CLK,
	output		    [23:0]		HDMI_TX_D,
	output		          		HDMI_TX_DE,
	output		          		HDMI_TX_HS,
	input 		          		HDMI_TX_INT,
	output		          		HDMI_TX_VS,

	// VGA
	output  [3:0] VGA_R,
	output  [3:0] VGA_G,
	output  [3:0] VGA_B,
	output        VGA_HS,
	output        VGA_VS
	
);



wire [31:0] status;
wire [1:0] buttons;

reg  direct = 1'b0;

// SELECT TYPE OF MEMORY ATTACHED
reg  [1:0] sdram_sz = 2'b01;       //0 - no memory board detected   1 - 32 MB  2 - 64 MB  3 - 128 MB



wire RESET = w_reset;

/*
wire joy1_up_i, joy1_down_i, joy1_left_i, joy1_right_i, joy1_p6_i, joy1_p9_i;
wire joy2_up_i, joy2_down_i, joy2_left_i, joy2_right_i, joy2_p6_i, joy2_p9_i;

joydecoder joystick_serial  (
    .clk          ( clock_50_i ), 	
    .joy_data     ( joy_data_i ),
    .joy_clk      ( joy_clock_o ),
    .joy_load     ( joy_load_o ),
	 .clock_locked ( locked ),

    .joy1up       ( joy1_up_i ),
    .joy1down     ( joy1_down_i ),
    .joy1left     ( joy1_left_i ),
    .joy1right    ( joy1_right_i ),
    .joy1fire1    ( joy1_p6_i ),
    .joy1fire2    ( joy1_p9_i ),

    .joy2up       ( joy2_up_i ),
    .joy2down     ( joy2_down_i ),
    .joy2left     ( joy2_left_i ),
    .joy2right    ( joy2_right_i ),
    .joy2fire1    ( joy2_p6_i ),
    .joy2fire2    ( joy2_p9_i )
); 
*/

///////////////////////////////////////////////////////////////////
wire clk_ram, locked;

wire [1:0] pll_locked_in;
wire pll_locked;
wire pll_areset;
wire pll_scanclk;
wire pll_scandata;
wire pll_scanclkena ;
wire pll_configupdate;
wire pll_scandataout;
wire pll_scandone;
wire [7:0]pll_rom_address;
wire pll_write_rom_ena;
wire pll_write_from_rom;
wire pll_reconfig_s;
wire pll_reconfig_busy;
wire pll_reconfig_reset;
reg [1:0]pll_reconfig_state = 2'b00;
integer pll_reconfig_timeout;
wire pll_rom_q;
	

pll pll
(
	
	.inclk0(clock_50_i),
	.areset(pll_areset | RESET),
	.c0(clk_ram),
	.c1(pll_clk),
	.locked(locked),
	
	.scanclk 		( pll_scanclk ),
	.scandata 		( pll_scandata ),
	.scanclkena 	( pll_scanclkena ),
	.configupdate 	( pll_configupdate ),
	.scandataout 	( pll_scandataout ),
	.scandone 		( pll_scandone )
	
);


	pll_reconfig pll_reconfig
	(
		.busy 					( pll_reconfig_busy ),
		.clock  					( clock_50_i ),
		.counter_param 		( 3'b000 ),
		.counter_type 			( 4'b0000 ),
		.data_in 				( 9'b000000000 ),
		.pll_areset 			( pll_areset ),
		.pll_areset_in  		( 0 ),
		.pll_configupdate 	( pll_configupdate),
		.pll_scanclk 			( pll_scanclk ),
		.pll_scanclkena 		( pll_scanclkena ),
		.pll_scandata 			( pll_scandata ),
		.pll_scandataout 		( pll_scandataout ),
      .pll_scandone		 	( pll_scandone ),
		.read_param			 	( 0 ),
      .reconfig 				( pll_reconfig_s ),
		.reset 					( pll_reconfig_reset ),
		.reset_rom_address 	( 0 ),
		.rom_address_out 		( pll_rom_address ),
		.rom_data_in 			( pll_rom_q ),
		.write_from_rom 		( pll_write_from_rom ),
		.write_param  			( 0 ),
      .write_rom_ena 		( pll_write_rom_ena )
	);
	

	wire q_reconfig_70, q_reconfig_80, q_reconfig_90, q_reconfig_100, q_reconfig_110, q_reconfig_120, q_reconfig_130, q_reconfig_140, q_reconfig_150, q_reconfig_160, q_reconfig_167;
	
	reconfig_70  reconfig_70  ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_70 ));
	reconfig_80  reconfig_80  ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_80 ));
	reconfig_90  reconfig_90  ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_90 ));
	reconfig_100 reconfig_100 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_100 ));
	reconfig_110 reconfig_110 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_110 ));
	reconfig_120 reconfig_120 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_120 ));
	reconfig_130 reconfig_130 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_130 ));
	reconfig_140 reconfig_140 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_140 ));
	reconfig_150 reconfig_150 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_150 ));
	reconfig_160 reconfig_160 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_160 ));
	reconfig_167 reconfig_167 ( .address ( pll_rom_address ), .clock ( clock_50_i ), .rden ( pll_write_rom_ena ), .q ( q_reconfig_167 ));

always @(*) 
begin
	case(pos)
		0: begin pll_rom_q <= q_reconfig_167; end
		1: begin pll_rom_q <= q_reconfig_160; end
		2: begin pll_rom_q <= q_reconfig_150; end
		3: begin pll_rom_q <= q_reconfig_140; end
		4: begin pll_rom_q <= q_reconfig_130; end
		5: begin pll_rom_q <= q_reconfig_120; end
		6: begin pll_rom_q <= q_reconfig_110; end
		7: begin pll_rom_q <= q_reconfig_100; end
		8: begin pll_rom_q <= q_reconfig_90;  end
		9: begin pll_rom_q <= q_reconfig_80;  end
	  10: begin pll_rom_q <= q_reconfig_70;  end
	endcase
end		

	
reg recfg = 0;

// Phases here are empirically adjusted based on 167MHz synthesized core 
// so arn't reliable for fixed frequency cores.
wire [31:0] cfg_param[44] =
'{ //      M         K          C
	'h167, 'h00808, 'hB33332DD, 'h20302,
	'h160, 'h00808, 'h00000001, 'h20302,
	'h150, 'h20807, 'h00000001, 'h20302,
	'h140, 'h00707, 'h00000001, 'h20302,
	'h130, 'h00505, 'h66666611, 'h00202,
	'h120, 'h00707, 'h66666611, 'h00303,
	'h110, 'h20706, 'h333332DD, 'h00303,
	'h100, 'h00404, 'h00000001, 'h00202,
	 'h90, 'h00707, 'h66666666, 'h00404,
	 'h80, 'h00707, 'h66666666, 'h20504,
	 'h70, 'h00707, 'h00000001, 'h00505
};

reg   [3:0] pos  = 7;
reg  [15:0] mins = 0;
reg  [15:0] secs = 0;
reg         auto = 0;

reg  [10:0] ps2_key;

reg btn_rst, old_btn_rst;
reg btn_up, old_btn_up;
reg btn_down, old_btn_down;
reg btn_auto, old_btn_auto;


always @(posedge clock_50_i) begin
	reg  [7:0] state = 0;
	integer    min = 0, sec = 0;
	reg        old_stb = 0;

	pll_write_from_rom <= 0;
	pll_reconfig_s <= 0;
	pll_reconfig_reset <= 0;





			case(pll_reconfig_state)
	
				0: begin
						if (recfg)
						begin
							pll_write_from_rom <= 1;
							pll_reconfig_state <= 1;
						end
					end

		
				1: begin
						pll_reconfig_state <= 2;
					end

			
				2: begin
				
						if (pll_reconfig_busy == 0)
						begin	
							pll_reconfig_s <= 1;
							pll_reconfig_state <= 3;
							pll_reconfig_timeout <= 1000;
						end;
						
					end

		
				3: begin
				
						pll_reconfig_timeout <= pll_reconfig_timeout - 1;
						
						if (pll_reconfig_timeout == 1) 
						begin
							pll_reconfig_reset <= 1; // sometimes pll reconfig stuck in busy state
							pll_reconfig_state <= 0;
							recfg <= 0;
						end
						
						if (pll_reconfig_s == 0 && pll_reconfig_busy == 0)
						begin
							pll_reconfig_state <= 0;
							recfg <= 0;
						end
						
					end


			endcase
	


	if(recfg) begin
		{min, mins} <= 0;
		{sec, secs} <= 0;
	end else begin
		min <= min + 1;
		if(min == 2999999999) begin
			min <= 0;
			if(mins[3:0]<9) mins[3:0] <= mins[3:0] + 1'd1;
			else begin
				mins[3:0] <= 0;
				if(mins[7:4]<9) mins[7:4] <= mins[7:4] + 1'd1;
				else begin
					mins[7:4] <= 0;
					if(mins[11:8]<9) mins[11:8] <= mins[11:8] + 1'd1;
					else begin
						mins[11:8] <= 0;
						if(mins[15:12]<9) mins[15:12] <= mins[15:12] + 1'd1;
						else mins[15:12] <= 0;
					end
				end
			end
		end
		sec <= sec + 1;
		if(sec == 4999999) begin
			sec <= 0;
			secs <= secs + 1'd1;
		end
	end
	
	old_btn_rst <= btn_rst;
	old_btn_up <= btn_up;
	old_btn_down <= btn_down;
	old_btn_auto <= btn_auto;
		
		//(pos 0 = 167)
		
	if(old_btn_rst == 0 && btn_rst == 1) 
	begin
	//	direct <= ~direct;
	end
	
		
	if(old_btn_up == 0 && btn_up == 1 && pos > 0) 
	begin
		state <= 0;
		recfg <= 1;
		pos <= pos - 1'd1;
		auto <= 0;
	end
			
	if(old_btn_down == 0 && btn_down == 1 && pos < 10) 
	begin
		state <= 0;
		recfg <= 1;
		pos <= pos + 1'd1;
		auto <= 0;
	end
			
	if(old_btn_auto == 0 && btn_auto == 1 && auto == 1) 
	begin
	state <= 0;
		recfg <= 1;
		auto <= 0;
	end
			
	if(old_btn_auto == 0 && btn_auto == 1 && auto == 0) 
	begin
		state <= 0;
		recfg <= 1;
		pos <= 0;
		auto <= 1;
	end

	if(auto && (failcount && passcount) && !recfg && pos < 10) 
	begin
		recfg <= 1;
		pos <= pos + 1'd1;
	end
	
	if(status[0] ) 
	begin
		recfg <= 1;
		pos <= 0;
		auto <= 1;
	end
end


///////////////////////////////////////////////////////////////////
assign SDRAM_CKE = 1;

reg reset = 0;
always @(posedge clk_ram) begin
	integer timeout;

	if(timeout) timeout <= timeout - 1;
	reset <= |timeout;

	if((recfg || ~locked) && (timeout < 1000000)) timeout <= 1000000;

	if(RESET) timeout <= 100000000;
end

wire module_clk, pll_clk;

wire [31:0] passcount, failcount;
tester my_memtst
(
	.clk(clk_ram),
	.rst_n(~reset),
	.sz(sdram_sz),
	.passcount(passcount),
	.failcount(failcount),
	.DRAM_CLK(SDRAM_CLK),
	.DRAM_DQ(SDRAM_DQ),
	.DRAM_ADDR(SDRAM_A),
	.DRAM_LDQM(SDRAM_DQML),
	.DRAM_UDQM(SDRAM_DQMH),
	.DRAM_WE_N(SDRAM_nWE),
	.DRAM_CS_N(SDRAM_nCS),
	.DRAM_RAS_N(SDRAM_nRAS),
	.DRAM_CAS_N(SDRAM_nCAS),
	.DRAM_BA_0(SDRAM_BA[0]),
	.DRAM_BA_1(SDRAM_BA[1])
);

///////////////////////////////////////////////////////////////////
//HDMI I2C	
I2C_HDMI_Config u_I2C_HDMI_Config (
	.iCLK(clock_50_i),
	.iRST_N(~RESET),
	.I2C_SCLK(HDMI_I2C_SCL),
	.I2C_SDAT(HDMI_I2C_SDA),
	.HDMI_TX_INT(HDMI_TX_INT)
	);

	assign HDMI_TX_DE = VGA_DE;
	assign HDMI_TX_HS = hs;
	assign HDMI_TX_VS = vs;	
	assign HDMI_TX_CLK = videoclk;
	assign HDMI_TX_D[23:16] = {8{r}};
	assign HDMI_TX_D[15:8] = {8{g}};
	assign HDMI_TX_D[7:0] = {8{b}};

///////////////////////////////////////////////////////////////////
// VGA VIDEO

wire videoclk;

vid_pll vid_pll
(
	.inclk0(clock_50_i),
	.c0(videoclk)
);

//assign CLK_VIDEO = videoclk;
//assign CE_PIXEL  = 1;

wire hs, vs, VGA_DE;
wire [1:0] b, r, g;

vgaout showrez
(
	.clk(videoclk),
	.rez1({(direct)?4'd13:4'd1, passcount[27:0]}),
	.rez2(failcount),
	.bg(6'b000001),
	.freq(16'hF000 | cfg_param[{pos, 2'd0}][11:0]),
	.elapsed(mins),
	.mark(8'h80 >> {~auto, secs[2:0]}),
	.hs(hs),
	.vs(vs),
	.de(VGA_DE),
	.b(b),
	.r(r),
	.g(g)
);

assign VGA_HS = ~hs;
assign VGA_VS = ~vs;

assign VGA_B  = {4{b}};
assign VGA_R  = {4{r}};
assign VGA_G  = {4{g}};

///////////////////////////////////////////////////////////////////

// delgrom keyboard and joysticks
wire [12:0] JoyPCFRLDU;
wire w_reset;

wire m_up     = JoyPCFRLDU[0] | ~KEY[0];   // | ~joy1_up_i;		//arriba
wire m_down   = JoyPCFRLDU[1] | ~KEY[1];   // | ~joy1_down_i;	//abajo
wire m_auto  =  JoyPCFRLDU[5] | ~SW[1];    // | ~joy1_p6_i;		//a
wire m_reset  =  w_reset;						//escape

debounce # ( .counter_size (10)) debounce1 ( .clk_i   (clock_50_i),   .button_i (m_reset), .result_o  (btn_rst)); 
debounce # ( .counter_size (10)) debounce2 ( .clk_i   (clock_50_i),   .button_i (m_up),   .result_o  (btn_up)); 
debounce # ( .counter_size (10)) debounce3 ( .clk_i   (clock_50_i),   .button_i (m_down), .result_o  (btn_down)); 
debounce # ( .counter_size (10)) debounce4 ( .clk_i   (clock_50_i),   .button_i (m_auto), .result_o  (btn_auto)); 

wire kbd_intr;
wire [7:0] kbd_scancode;
wire [7:0] keys_s;

//get scancode from keyboard
io_ps2_keyboard keyboard 
 (
  .clk       ( clock_50_i ),
  .kbd_clk   ( ps2_clk_io ),
  .kbd_dat   ( ps2_data_io ),
  .interrupt ( kbd_intr ),
  .scancode  ( kbd_scancode )
);

//translate scancode to joystick
kbd_joystick k_joystick
(
  .clk         	( clock_50_i ),
  .kbdint      	( kbd_intr ),
  .kbdscancode 	( kbd_scancode ), 
  .JoyPCFRLDU     ( JoyPCFRLDU ),
  .osd_o	  ( keys_s ),
  .reset          (w_reset)
);


endmodule
